1,small
6,size 2
7,size 3
8,size 4
9,size 5
